module PATTERN_GENERATOR_HANDLE
(
	input					CLK_100MHz,
	input					nRESET,
	input		[7:1]		ADDRESS,
	inout		[15:0]	DATA,
	input					nCS,
	input					nRE,
	input					nWE,
	
	input					REF_CLK,
	input					SYNC,
	//input					PATTERN_ON,
	output 				OUTPUT_nON,
	output	[23:0]	LEVEL_SEL,
	output				INTERRUPT,
	output				DAC_LOAD_CONTROL
);

parameter	BASE_ADDRESS				=		7'd50,
				STATUS_OFFSET				=		7'd0,
				CONTROL_OFFSET				=		7'd1,
				VTOTAL_L_OFFSET			=		7'd2,
				VTOTAL_H_OFFSET			=		7'd3,
				INVERSION_L_OFFSET		=		7'd4,
				INVERSION_H_OFFSET		=		7'd5,
				SET_L_OFFSET				=		7'd6,
				SET_H_OFFSET				=		7'd7,
				DELAY_VALUE_L				=		7'd8,
				DELAY_VALUE_H				=		7'd9,
				WIDTH_VALUE_L				=		7'd10,
				WIDTH_VALUE_H				=		7'd11,
				PERIOD_VALUE_L				=		7'd12,
				PERIOD_VALUE_H				=		7'd13,
				START_VALUE_L				=		7'd14,
				START_VALUE_H				=		7'd15,
				END_VALUE_L					=		7'd16,
				END_VALUE_H					=		7'd17,
				OUTPUT_DELAY_L				=		7'd18,
				OUTPUT_DELAY_H				=		7'd19;
				
/*
STATUS
bit 1~15 Reseved
bit 1 analog Mux Enbale
bit 0 pattern on
*/
reg		[15:0]			REG_STATUS;
/*
CONTROL
bit 8~15 Reseved
bit 7 VR_RGB_ON
bit 6 Force Pattern_ON
bit 5 SYNC
bit 4 INTERRUPT_ON
bit 3 TIMING_CHANGE
buf 2 INVERSION_CHANGE
bit 1 PARRTERN_CHANGE for DAC_LOAD
bit 0 PATTERN_ON for Analog MUX nENABLE
*/
reg		[15:0]			REG_CONTROL;
reg		[15:0]			REG_VTOTAL_L;
reg		[15:0]			REG_VTOTAL_H;
wire		[31:0]			WIRE_VTOTAL;
assign WIRE_VTOTAL = {REG_VTOTAL_H, REG_VTOTAL_L};
reg		[31:0]			BUF_VTOTAL;
reg		[15:0]			REG_INVERSION_L;
reg		[15:0]			REG_INVERSION_H;
reg		[31:0]			BUF_INVERSION;
reg		[15:0]			REG_SET_L;
reg		[15:0]			REG_SET_H;
wire		[31:0]			WIRE_SET;
assign	WIRE_SET = {REG_SET_H, REG_SET_L};
reg		[15:0]			REG_DELAY_VALUE_L;
reg		[15:0]			REG_DELAY_VALUE_H;
wire		[31:0]			WIRE_DELAY;
assign	WIRE_DELAY = {REG_DELAY_VALUE_H, REG_DELAY_VALUE_L};
reg		[15:0]			REG_WIDTH_VALUE_L;
reg		[15:0]			REG_WIDTH_VALUE_H;
wire		[31:0]			WIRE_WIDTH;
assign	WIRE_WIDTH = {REG_WIDTH_VALUE_H, REG_WIDTH_VALUE_L};
reg		[15:0]			REG_PERIOD_VALUE_L;
reg		[15:0]			REG_PERIOD_VALUE_H;
wire		[31:0]			WIRE_PERIOD;
assign	WIRE_PERIOD = {REG_PERIOD_VALUE_H, REG_PERIOD_VALUE_L};
reg		[15:0]			REG_START_VALUE_L;
reg		[15:0]			REG_START_VALUE_H;
wire		[31:0]			WIRE_START;
assign	WIRE_START = {REG_START_VALUE_H, REG_START_VALUE_L};
reg		[15:0]			REG_END_VALUE_L;
reg		[15:0]			REG_END_VALUE_H;
wire		[31:0]			WIRE_END;
assign	WIRE_END = {REG_END_VALUE_H, REG_END_VALUE_L};
reg		[15:0]			REG_OUTPUT_DELAY_L;
reg		[15:0]			REG_OUTPUT_DELAY_H;
wire		[31:0]			WIRE_OUTPUT_DELAY;
assign	WIRE_OUTPUT_DELAY = {REG_OUTPUT_DELAY_H, REG_OUTPUT_DELAY_L};

always @ (posedge CLK_100MHz) begin
	if(!nRESET) begin
		REG_STATUS <= 16'b0000000000000000;
		REG_CONTROL <= 16'b0000000000110000;
		REG_SET_L <= 16'b0000000000000000;
		REG_SET_H <= 16'b0000000000000000;
		REG_DELAY_VALUE_L <= 16'b0000000000000000;
		REG_DELAY_VALUE_H <= 16'b0000000000000000;
		REG_WIDTH_VALUE_L <= 16'b0000000000000000;
		REG_WIDTH_VALUE_H <= 16'b0000000000000000;
		REG_PERIOD_VALUE_L <= 16'b0000000000000000;
		REG_PERIOD_VALUE_H <= 16'b0000000000000000;
		REG_START_VALUE_L <= 16'b0000000000000000;
		REG_START_VALUE_H <= 16'b0000000000000000;
		REG_END_VALUE_L <= 16'b0000000000000000;
		REG_END_VALUE_H <= 16'b0000000000000000;
		REG_OUTPUT_DELAY_L <= 16'd0;
		REG_OUTPUT_DELAY_H <= 16'd0;
	end
	else begin
		if((!nCS) && (!nWE)) begin
			if			(ADDRESS == (BASE_ADDRESS + CONTROL_OFFSET))					REG_CONTROL					<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + VTOTAL_L_OFFSET))				REG_VTOTAL_L				<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + VTOTAL_H_OFFSET))				REG_VTOTAL_H				<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + INVERSION_L_OFFSET))			REG_INVERSION_L			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + INVERSION_H_OFFSET))			REG_INVERSION_H			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + SET_L_OFFSET))					REG_SET_L					<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + SET_H_OFFSET))					REG_SET_H					<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DELAY_VALUE_L))					REG_DELAY_VALUE_L			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DELAY_VALUE_H))					REG_DELAY_VALUE_H			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + WIDTH_VALUE_L))					REG_WIDTH_VALUE_L			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + WIDTH_VALUE_H))					REG_WIDTH_VALUE_H			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + PERIOD_VALUE_L))					REG_PERIOD_VALUE_L		<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + PERIOD_VALUE_H))					REG_PERIOD_VALUE_H		<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + START_VALUE_L))					REG_START_VALUE_L			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + START_VALUE_H))					REG_START_VALUE_H			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + END_VALUE_L))						REG_END_VALUE_L			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + END_VALUE_H))						REG_END_VALUE_H			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + OUTPUT_DELAY_L))					REG_OUTPUT_DELAY_L		<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + OUTPUT_DELAY_H))					REG_OUTPUT_DELAY_H		<=		DATA;
		end
		if(REG_DAC_LOAD_DONE == 10'b1111111111) REG_CONTROL[1] <= 1'd0;
		if(WIRE_SETTING_DONE[0] == 1'b1) REG_CONTROL[2] <= 1'd0;
		if(WIRE_SETTING_DONE[1] == 1'b1) REG_CONTROL[3] <= 1'd0;
		if(REG_VR_RGB_OPERATION == 1'b1) REG_CONTROL[7] <= 1'd0;
		//REG_STATUS[0] <= ~PATTERN_ON;
		REG_STATUS[0] <= REG_CONTROL[0];
		REG_STATUS[1] <= ~REG_OUTPUT_nON;
	end
end

wire		[15:0]		READ_DATA;
assign	DATA			=		(!nCS && !nRE) ? READ_DATA : 16'bzzzzzzzzzzzzzzzz;
assign	READ_DATA	=		(ADDRESS == (BASE_ADDRESS + STATUS_OFFSET))					?		REG_STATUS :
									(ADDRESS == (BASE_ADDRESS + CONTROL_OFFSET))					?		REG_CONTROL :
									(ADDRESS == (BASE_ADDRESS + VTOTAL_L_OFFSET))				?		REG_VTOTAL_L :
									(ADDRESS == (BASE_ADDRESS + VTOTAL_H_OFFSET))				?		REG_VTOTAL_H :
									(ADDRESS == (BASE_ADDRESS + INVERSION_L_OFFSET))			?		REG_INVERSION_L :
									(ADDRESS == (BASE_ADDRESS + INVERSION_H_OFFSET))			?		REG_INVERSION_H :
									(ADDRESS == (BASE_ADDRESS + SET_L_OFFSET))					?		REG_SET_L :
									(ADDRESS == (BASE_ADDRESS + SET_H_OFFSET))					?		REG_SET_H :
									(ADDRESS == (BASE_ADDRESS + DELAY_VALUE_L))					?		REG_DELAY_VALUE_L :
									(ADDRESS == (BASE_ADDRESS + DELAY_VALUE_H))					?		REG_DELAY_VALUE_H :
									(ADDRESS == (BASE_ADDRESS + WIDTH_VALUE_L))					?		REG_WIDTH_VALUE_L :
									(ADDRESS == (BASE_ADDRESS + WIDTH_VALUE_H))					?		REG_WIDTH_VALUE_H :
									(ADDRESS == (BASE_ADDRESS + PERIOD_VALUE_L))					?		REG_PERIOD_VALUE_L :
									(ADDRESS == (BASE_ADDRESS + PERIOD_VALUE_H))					?		REG_PERIOD_VALUE_H :
									(ADDRESS == (BASE_ADDRESS + START_VALUE_L))					?		REG_START_VALUE_L :
									(ADDRESS == (BASE_ADDRESS + START_VALUE_H))					?		REG_START_VALUE_H :
									(ADDRESS == (BASE_ADDRESS + END_VALUE_L))						?		REG_END_VALUE_L :
									(ADDRESS == (BASE_ADDRESS + END_VALUE_H))						?		REG_END_VALUE_L :
									(ADDRESS == (BASE_ADDRESS + OUTPUT_DELAY_L))					?		REG_OUTPUT_DELAY_L :
									(ADDRESS == (BASE_ADDRESS + OUTPUT_DELAY_H))					?		REG_OUTPUT_DELAY_H : 16'bzzzzzzzzzzzzzzzz;

assign INTERRUPT = REG_CONTROL[4];
wire							WIRE_VSYNC;
wire							WIRE_SYNC;
assign WIRE_SYNC = REG_CONTROL[5] & SYNC;

//reg REG_PATTERN_ON;
reg [1:0] REG_VSYNC_DETECT;
always @ (posedge REF_CLK) begin
	if(!nRESET) begin
		//REG_PATTERN_ON <= 1'd0;
		REG_VSYNC_DETECT <= 2'b11;
	end
	else begin
		//if(!PATTERN_ON) REG_PATTERN_ON <= 1'd1;
		//else REG_PATTERN_ON <= 1'd0;
		REG_VSYNC_DETECT <= {REG_VSYNC_DETECT[0], WIRE_VSYNC};
	end
end

reg REG_OUTPUT_nON;
reg [1:0] REG_OUTPUT_nON_DELAY;
assign OUTPUT_nON = REG_OUTPUT_nON_DELAY[1];
reg REG_DAC_LOAD_CONTROL;
reg [1:0] REG_DAC_LOAD_CONTROL_DELAY;
assign DAC_LOAD_CONTROL = REG_DAC_LOAD_CONTROL_DELAY[1];
reg [9:0] REG_DAC_LOAD_DONE;
reg [1:0] REG_SETTING_CHANGE;
wire [23:0] WIRE_SETTING_INVESION_DONE_ARRAY;
wire [23:0] WIRE_SETTING_TIMING_DONE_ARRAY;
wire	[1:0] WIRE_SETTING_DONE;
assign WIRE_SETTING_DONE[0] = WIRE_SETTING_INVESION_DONE_ARRAY[0] & WIRE_SETTING_INVESION_DONE_ARRAY[1] & WIRE_SETTING_INVESION_DONE_ARRAY[2] & WIRE_SETTING_INVESION_DONE_ARRAY[3]
									& WIRE_SETTING_INVESION_DONE_ARRAY[4] & WIRE_SETTING_INVESION_DONE_ARRAY[5] & WIRE_SETTING_INVESION_DONE_ARRAY[6] & WIRE_SETTING_INVESION_DONE_ARRAY[7]
									& WIRE_SETTING_INVESION_DONE_ARRAY[8] & WIRE_SETTING_INVESION_DONE_ARRAY[9] & WIRE_SETTING_INVESION_DONE_ARRAY[10] & WIRE_SETTING_INVESION_DONE_ARRAY[11]
									& WIRE_SETTING_INVESION_DONE_ARRAY[12] & WIRE_SETTING_INVESION_DONE_ARRAY[13] & WIRE_SETTING_INVESION_DONE_ARRAY[14] & WIRE_SETTING_INVESION_DONE_ARRAY[15]
									& WIRE_SETTING_INVESION_DONE_ARRAY[16] & WIRE_SETTING_INVESION_DONE_ARRAY[17] & WIRE_SETTING_INVESION_DONE_ARRAY[18] & WIRE_SETTING_INVESION_DONE_ARRAY[19]
									& WIRE_SETTING_INVESION_DONE_ARRAY[20] & WIRE_SETTING_INVESION_DONE_ARRAY[21] & WIRE_SETTING_INVESION_DONE_ARRAY[22] & WIRE_SETTING_INVESION_DONE_ARRAY[23];
assign WIRE_SETTING_DONE[1] = WIRE_SETTING_TIMING_DONE_ARRAY[0] & WIRE_SETTING_TIMING_DONE_ARRAY[1] & WIRE_SETTING_TIMING_DONE_ARRAY[2] & WIRE_SETTING_TIMING_DONE_ARRAY[3]
									& WIRE_SETTING_TIMING_DONE_ARRAY[4] & WIRE_SETTING_TIMING_DONE_ARRAY[5] & WIRE_SETTING_TIMING_DONE_ARRAY[6] & WIRE_SETTING_TIMING_DONE_ARRAY[7]
									& WIRE_SETTING_TIMING_DONE_ARRAY[8] & WIRE_SETTING_TIMING_DONE_ARRAY[9] & WIRE_SETTING_TIMING_DONE_ARRAY[10] & WIRE_SETTING_TIMING_DONE_ARRAY[11]
									& WIRE_SETTING_TIMING_DONE_ARRAY[12] & WIRE_SETTING_TIMING_DONE_ARRAY[13] & WIRE_SETTING_TIMING_DONE_ARRAY[14] & WIRE_SETTING_TIMING_DONE_ARRAY[15]
									& WIRE_SETTING_TIMING_DONE_ARRAY[16] & WIRE_SETTING_TIMING_DONE_ARRAY[17] & WIRE_SETTING_TIMING_DONE_ARRAY[18] & WIRE_SETTING_TIMING_DONE_ARRAY[19]
									& WIRE_SETTING_TIMING_DONE_ARRAY[20] & WIRE_SETTING_TIMING_DONE_ARRAY[21] & WIRE_SETTING_TIMING_DONE_ARRAY[22] & WIRE_SETTING_TIMING_DONE_ARRAY[23];

reg REG_SYNC_OPERATION;
reg REG_VR_RGB_OPERATION;

reg [1:0] REG_WIRE_SYNC_NEG_CATCH;
always @ (negedge CLK_100MHz) begin
	if(!nRESET) begin
		REG_WIRE_SYNC_NEG_CATCH <= 2'b00;
	end
	else begin
		REG_WIRE_SYNC_NEG_CATCH <= {REG_WIRE_SYNC_NEG_CATCH[0], WIRE_SYNC};
	end
end

always @ (posedge CLK_100MHz) begin
	if(!nRESET) begin
		REG_OUTPUT_nON <= 1'd1;
		REG_DAC_LOAD_CONTROL <= 1'b1;
		REG_DAC_LOAD_DONE <= 10'b0000000000;
		REG_SETTING_CHANGE <= 2'b00;
		BUF_INVERSION <= 32'd0;
		BUF_VTOTAL <= 32'd10;
		REG_SYNC_OPERATION <= 1'd0;
		REG_VR_RGB_OPERATION <= 1'd0;
	end
	else begin
		if((REG_WIRE_SYNC_NEG_CATCH[1] == 1'b1) && (REG_WIRE_SYNC_NEG_CATCH[0] == 1'b0)) REG_SYNC_OPERATION <= 1'd1;
		else begin
			if((REG_SYNC_OPERATION) || (REG_CONTROL[7]))begin
				if((REG_VSYNC_DETECT[1] == 1'd0) && (REG_VSYNC_DETECT[0] == 1'd1)) begin
					REG_SYNC_OPERATION <= 1'd0;
					REG_VR_RGB_OPERATION <= 1'd1;
					//if((REG_PATTERN_ON && REG_CONTROL[0]) || (REG_CONTROL[6])) REG_OUTPUT_nON <= 1'd0;
					if((REG_CONTROL[0]) || (REG_CONTROL[6])) REG_OUTPUT_nON <= 1'd0;
					else REG_OUTPUT_nON <= 1'd1;
					if(REG_CONTROL[1]) REG_DAC_LOAD_CONTROL <= 1'd0;
					if(REG_CONTROL[2]) begin
						BUF_INVERSION <= {REG_INVERSION_H, REG_INVERSION_L};
						REG_SETTING_CHANGE[0] <= 1'd1;
					end
				end
				if(REG_CONTROL[3]) begin
					REG_SETTING_CHANGE[1] <= 1'd1;
					if(WIRE_VTOTAL >= 32'd10) BUF_VTOTAL <= {REG_VTOTAL_H, REG_VTOTAL_L};
					else BUF_VTOTAL <= 32'd10;
				end
			end
			else begin
				if(!REG_DAC_LOAD_CONTROL) REG_DAC_LOAD_DONE <= {REG_DAC_LOAD_DONE[8:0], 1'd1};
				if(!REG_CONTROL[1]) begin
					REG_DAC_LOAD_CONTROL <= 1'd1;
					REG_DAC_LOAD_DONE <= 10'b0000000000;
				end
				if(!REG_CONTROL[2]) REG_SETTING_CHANGE[0] <= 1'd0;
				if(!REG_CONTROL[3]) REG_SETTING_CHANGE[1] <= 1'd0;
				if(!REG_CONTROL[7]) REG_VR_RGB_OPERATION <= 1'd0;
			end
		end
	end
end

always @ (posedge REF_CLK) begin //OUTPUT_nON, DAC_LOAD : 2Clock Delay
	if(!nRESET) begin
		REG_DAC_LOAD_CONTROL_DELAY <= 2'b11;
		REG_OUTPUT_nON_DELAY <= 2'b11;
	end
	else begin
		REG_DAC_LOAD_CONTROL_DELAY <= {REG_DAC_LOAD_CONTROL_DELAY[0], REG_DAC_LOAD_CONTROL};
		REG_OUTPUT_nON_DELAY <= {REG_OUTPUT_nON_DELAY[0], REG_OUTPUT_nON};
	end
end

VSYNC_GENERATOR VSYNC_GENERATOR_inst
(
	.nRESET(nRESET) ,	// input  nRESET_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.SYNC(WIRE_SYNC) ,	// input  SYNC_sig
	.VTOTAL(BUF_VTOTAL) ,	// input [31:0] VTOTAL_sig
	.DELAY(WIRE_OUTPUT_DELAY) ,	// input [31:0] DELAY_sig
	.VSYNC(WIRE_VSYNC) 	// output  VSYNC_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst0
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[0]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[0], WIRE_SETTING_INVESION_DONE_ARRAY[0]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[0]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[0]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst1
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[1]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[1], WIRE_SETTING_INVESION_DONE_ARRAY[1]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[1]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[1]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst2
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[2]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[2], WIRE_SETTING_INVESION_DONE_ARRAY[2]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[2]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[2]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst3
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[3]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[3], WIRE_SETTING_INVESION_DONE_ARRAY[3]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[3]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[3]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst4
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[4]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[4], WIRE_SETTING_INVESION_DONE_ARRAY[4]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[4]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[4]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst5
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[5]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[5], WIRE_SETTING_INVESION_DONE_ARRAY[5]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[5]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[5]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst6
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[6]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[6], WIRE_SETTING_INVESION_DONE_ARRAY[6]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[6]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[6]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst7
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[7]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[7], WIRE_SETTING_INVESION_DONE_ARRAY[7]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[7]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[7]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst8
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[8]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[8], WIRE_SETTING_INVESION_DONE_ARRAY[8]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[8]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[8]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst9
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[9]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[9], WIRE_SETTING_INVESION_DONE_ARRAY[9]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[9]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[9]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst10
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[10]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[10], WIRE_SETTING_INVESION_DONE_ARRAY[10]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[10]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[10]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst11
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[11]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[11], WIRE_SETTING_INVESION_DONE_ARRAY[11]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[11]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[11]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst12
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[12]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[12], WIRE_SETTING_INVESION_DONE_ARRAY[12]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[12]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[12]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst13
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[13]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[13], WIRE_SETTING_INVESION_DONE_ARRAY[13]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[13]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[13]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst14
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[14]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[14], WIRE_SETTING_INVESION_DONE_ARRAY[14]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[14]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[14]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst15
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[15]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[15], WIRE_SETTING_INVESION_DONE_ARRAY[15]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[15]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[15]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst16
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[16]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[16], WIRE_SETTING_INVESION_DONE_ARRAY[16]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[16]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[16]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst17
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[17]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[17], WIRE_SETTING_INVESION_DONE_ARRAY[17]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[17]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[17]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst18
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[18]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[18], WIRE_SETTING_INVESION_DONE_ARRAY[18]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[18]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[18]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst19
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[19]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[19], WIRE_SETTING_INVESION_DONE_ARRAY[19]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[19]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[19]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst20
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[20]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[20], WIRE_SETTING_INVESION_DONE_ARRAY[20]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[20]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[20]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst21
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[21]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[21], WIRE_SETTING_INVESION_DONE_ARRAY[21]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[21]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[21]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst22
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[22]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[22], WIRE_SETTING_INVESION_DONE_ARRAY[22]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[22]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[22]) 	// output  LEVEL_SEL_sig
);

TIMING_GENERATOR TIMING_GENERATOR_inst23
(
	//.OUT_CLK(CLK_100MHz) , // input OUT_CLK_sig
	.REF_CLK(REF_CLK) ,	// input  REF_CLK_sig
	.nRESET(nRESET) ,	// input  nRESET_sig
	.SET(WIRE_SET[23]) ,	// input  SET_sig
	.DELAY(WIRE_DELAY) ,	// input [31:0] DELAY_sig
	.WIDTH(WIRE_WIDTH) ,	// input [31:0] WIDTH_sig
	.PERIOD(WIRE_PERIOD) ,	// input [31:0] PERIOD_sig
	.START(WIRE_START) ,	// input [31:0] START_sig
	.END(WIRE_END) ,	// input [31:0] END_sig
	.SETTING_EN(REG_SETTING_CHANGE) ,	// input SETTING_EN_sig
	.SETTING_DONE({WIRE_SETTING_TIMING_DONE_ARRAY[23], WIRE_SETTING_INVESION_DONE_ARRAY[23]}) ,	// input SETTING_DONE_sig
	.VSYNC(WIRE_VSYNC) ,	// input  VSYNC_sig
	.INVERSION_EN(BUF_INVERSION[23]) ,	// input  INVERSION_EN_sig
	.LEVEL_SEL(LEVEL_SEL[23]) 	// output  LEVEL_SEL_sig
);

endmodule
