module DAC_HANDLE
(
	input					CLK_100MHz,
	input					nRESET,
	input		[7:1]		ADDRESS,
	inout		[15:0]	DATA,
	input					nCS,
	input					nRE,
	input					nWE,
	
	input					DAC_REF_CLK,
	output	[4:0]		DAC_SCLK,
	output	[4:0]		DAC_nCS,
	output				DAC_SDI,
	output				DAC_nRST,
	output				DAC_nLOAD,
	
	input					EXTERNAL_DAC_nLOAD
);

parameter	BASE_ADDRESS				=		7'd0,

				DAC_STATUS_OFFSET			=		7'd0,
				DAC_CONTROL_OFFSET		=		7'd1,
				DAC0_OUTPUT0_OFFSET		=		7'd2,
				DAC0_OUTPUT1_OFFSET		=		7'd3,
				DAC0_OUTPUT2_OFFSET		=		7'd4,
				DAC0_OUTPUT3_OFFSET		=		7'd5,
				DAC1_OUTPUT0_OFFSET		=		7'd6,
				DAC1_OUTPUT1_OFFSET		=		7'd7,
				DAC1_OUTPUT2_OFFSET		=		7'd8,
				DAC1_OUTPUT3_OFFSET		=		7'd9,
				DAC2_OUTPUT0_OFFSET		=		7'd10,
				DAC2_OUTPUT1_OFFSET		=		7'd11,
				DAC2_OUTPUT2_OFFSET		=		7'd12,
				DAC2_OUTPUT3_OFFSET		=		7'd13,
				DAC3_OUTPUT0_OFFSET		=		7'd14,
				DAC3_OUTPUT1_OFFSET		=		7'd15,
				DAC3_OUTPUT2_OFFSET		=		7'd16,
				DAC3_OUTPUT3_OFFSET		=		7'd17,
				DAC4_OUTPUT0_OFFSET		=		7'd18,
				DAC4_OUTPUT1_OFFSET		=		7'd19,
				DAC4_OUTPUT2_OFFSET		=		7'd20,
				DAC4_OUTPUT3_OFFSET		=		7'd21,
				DAC_SETCONTROL_OFFSET	=		7'd22,
				DAC_SETBUFFER0_OFFSET	=		7'd23,
				DAC_SETBUFFER1_OFFSET	=		7'd24;

/*
DAC_STATUS
bit 1~15 Reserved
bit 0 DAC_nREADY
*/
reg		[15:0]			REG_DAC_STATUS;
/*
DAC_CONTROL
bit 3~15 Reseved
bit 2 DAC_LD
bit 1 DAC_RST
bit 0 DAC_TX_START
*/
reg		[15:0]			REG_DAC_CONTROL;

reg		[15:0]			REG_DAC0_OUTPUT0;
reg		[15:0]			REG_DAC0_OUTPUT1;
reg		[15:0]			REG_DAC0_OUTPUT2;
reg		[15:0]			REG_DAC0_OUTPUT3;
reg		[15:0]			REG_DAC1_OUTPUT0;
reg		[15:0]			REG_DAC1_OUTPUT1;
reg		[15:0]			REG_DAC1_OUTPUT2;
reg		[15:0]			REG_DAC1_OUTPUT3;
reg		[15:0]			REG_DAC2_OUTPUT0;
reg		[15:0]			REG_DAC2_OUTPUT1;
reg		[15:0]			REG_DAC2_OUTPUT2;
reg		[15:0]			REG_DAC2_OUTPUT3;
reg		[15:0]			REG_DAC3_OUTPUT0;
reg		[15:0]			REG_DAC3_OUTPUT1;
reg		[15:0]			REG_DAC3_OUTPUT2;
reg		[15:0]			REG_DAC3_OUTPUT3;
reg		[15:0]			REG_DAC4_OUTPUT0;
reg		[15:0]			REG_DAC4_OUTPUT1;
reg		[15:0]			REG_DAC4_OUTPUT2;
reg		[15:0]			REG_DAC4_OUTPUT3;

/*
DAC_SETCONTROL default : b'0000000000000000 0x0000
bit 0~4 DAC_SET_START
*/
reg		[15:0]			REG_DAC_SETCONTROL;
reg		[15:0]			REG_DAC_SETBUFFER0;
reg		[15:0]			REG_DAC_SETBUFFER1;	

wire							WIRE_OUTPUT_DONE;
wire							WIRE_SET_DONE;
wire							WIRE_READY;

always @ (posedge CLK_100MHz) begin
	if(!nRESET) begin
		REG_DAC_STATUS			<=			16'b0000000000000001;
		REG_DAC_CONTROL		<=			16'b0000000000000000;
		REG_DAC_SETCONTROL	<=			16'b0000000000000000;
	end
	else begin
		if((!nCS) && (!nWE)) begin
			if			(ADDRESS == (BASE_ADDRESS + DAC_CONTROL_OFFSET))			REG_DAC_CONTROL			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC0_OUTPUT0_OFFSET))			REG_DAC0_OUTPUT0			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC0_OUTPUT1_OFFSET))			REG_DAC0_OUTPUT1			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC0_OUTPUT2_OFFSET))			REG_DAC0_OUTPUT2			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC0_OUTPUT3_OFFSET))			REG_DAC0_OUTPUT3			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC1_OUTPUT0_OFFSET))			REG_DAC1_OUTPUT0			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC1_OUTPUT1_OFFSET))			REG_DAC1_OUTPUT1			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC1_OUTPUT2_OFFSET))			REG_DAC1_OUTPUT2			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC1_OUTPUT3_OFFSET))			REG_DAC1_OUTPUT3			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC2_OUTPUT0_OFFSET))			REG_DAC2_OUTPUT0			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC2_OUTPUT1_OFFSET))			REG_DAC2_OUTPUT1			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC2_OUTPUT2_OFFSET))			REG_DAC2_OUTPUT2			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC2_OUTPUT3_OFFSET))			REG_DAC2_OUTPUT3			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC3_OUTPUT0_OFFSET))			REG_DAC3_OUTPUT0			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC3_OUTPUT1_OFFSET))			REG_DAC3_OUTPUT1			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC3_OUTPUT2_OFFSET))			REG_DAC3_OUTPUT2			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC3_OUTPUT3_OFFSET))			REG_DAC3_OUTPUT3			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC4_OUTPUT0_OFFSET))			REG_DAC4_OUTPUT0			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC4_OUTPUT1_OFFSET))			REG_DAC4_OUTPUT1			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC4_OUTPUT2_OFFSET))			REG_DAC4_OUTPUT2			<=		DATA;
			else if	(ADDRESS	== (BASE_ADDRESS + DAC4_OUTPUT3_OFFSET))			REG_DAC4_OUTPUT3			<=		DATA;
			else if	(ADDRESS == (BASE_ADDRESS + DAC_SETCONTROL_OFFSET))		REG_DAC_SETCONTROL		<=		DATA;
			else if	(ADDRESS == (BASE_ADDRESS + DAC_SETBUFFER0_OFFSET))		REG_DAC_SETBUFFER0		<=		DATA;
			else if	(ADDRESS == (BASE_ADDRESS + DAC_SETBUFFER1_OFFSET))		REG_DAC_SETBUFFER1		<=		DATA;
		end
		if(WIRE_OUTPUT_DONE) REG_DAC_CONTROL[0] <= 1'b0;
		if(INTERNAL_DAC_nRESET_DONE == 3'b111) REG_DAC_CONTROL[1] <= 1'b0;
		if(INTERNAL_DAC_nLOAD_DONE == 3'b111) REG_DAC_CONTROL[2] <= 1'b0;
		if(WIRE_SET_DONE) REG_DAC_SETCONTROL[4:0] <= 5'b00000;
		REG_DAC_STATUS[0] <= WIRE_READY;
	end
end

wire		[15:0]		READ_DATA;
assign	DATA			=		(!nCS && !nRE) ? READ_DATA : 16'bzzzzzzzzzzzzzzzz;
assign	READ_DATA	=		(ADDRESS == (BASE_ADDRESS + DAC_STATUS_OFFSET))			?		REG_DAC_STATUS :
									(ADDRESS == (BASE_ADDRESS + DAC_CONTROL_OFFSET))		?		REG_DAC_CONTROL :
									(ADDRESS == (BASE_ADDRESS + DAC0_OUTPUT0_OFFSET))		?		REG_DAC0_OUTPUT0 :
									(ADDRESS == (BASE_ADDRESS + DAC0_OUTPUT1_OFFSET))		?		REG_DAC0_OUTPUT1 :
									(ADDRESS == (BASE_ADDRESS + DAC0_OUTPUT2_OFFSET))		?		REG_DAC0_OUTPUT2 :
									(ADDRESS == (BASE_ADDRESS + DAC0_OUTPUT3_OFFSET))		?		REG_DAC0_OUTPUT3 :
									(ADDRESS == (BASE_ADDRESS + DAC1_OUTPUT0_OFFSET))		?		REG_DAC1_OUTPUT0 :
									(ADDRESS == (BASE_ADDRESS + DAC1_OUTPUT1_OFFSET))		?		REG_DAC1_OUTPUT1 :
									(ADDRESS == (BASE_ADDRESS + DAC1_OUTPUT2_OFFSET))		?		REG_DAC1_OUTPUT2 :
									(ADDRESS == (BASE_ADDRESS + DAC1_OUTPUT3_OFFSET))		?		REG_DAC1_OUTPUT3 :
									(ADDRESS == (BASE_ADDRESS + DAC2_OUTPUT0_OFFSET))		?		REG_DAC2_OUTPUT0 :
									(ADDRESS == (BASE_ADDRESS + DAC2_OUTPUT1_OFFSET))		?		REG_DAC2_OUTPUT1 :
									(ADDRESS == (BASE_ADDRESS + DAC2_OUTPUT2_OFFSET))		?		REG_DAC2_OUTPUT2 :
									(ADDRESS == (BASE_ADDRESS + DAC2_OUTPUT3_OFFSET))		?		REG_DAC2_OUTPUT3 :
									(ADDRESS == (BASE_ADDRESS + DAC3_OUTPUT0_OFFSET))		?		REG_DAC3_OUTPUT0 :
									(ADDRESS == (BASE_ADDRESS + DAC3_OUTPUT1_OFFSET))		?		REG_DAC3_OUTPUT1 :
									(ADDRESS == (BASE_ADDRESS + DAC3_OUTPUT2_OFFSET))		?		REG_DAC3_OUTPUT2 :
									(ADDRESS == (BASE_ADDRESS + DAC3_OUTPUT3_OFFSET))		?		REG_DAC3_OUTPUT3 :
									(ADDRESS == (BASE_ADDRESS + DAC4_OUTPUT0_OFFSET))		?		REG_DAC4_OUTPUT0 :
									(ADDRESS == (BASE_ADDRESS + DAC4_OUTPUT1_OFFSET))		?		REG_DAC4_OUTPUT1 :
									(ADDRESS == (BASE_ADDRESS + DAC4_OUTPUT2_OFFSET))		?		REG_DAC4_OUTPUT2 :
									(ADDRESS == (BASE_ADDRESS + DAC4_OUTPUT3_OFFSET))		?		REG_DAC4_OUTPUT3 :
									(ADDRESS == (BASE_ADDRESS + DAC_SETCONTROL_OFFSET))	?		REG_DAC_SETCONTROL :
									(ADDRESS == (BASE_ADDRESS + DAC_SETBUFFER0_OFFSET))	?		REG_DAC_SETBUFFER0 :
									(ADDRESS == (BASE_ADDRESS + DAC_SETBUFFER1_OFFSET))	?		REG_DAC_SETBUFFER1 : 16'bzzzzzzzzzzzzzzzz;

reg INTERNAL_DAC_nRESET;
reg [2:0] INTERNAL_DAC_nRESET_DONE;
reg INTERNAL_DAC_nLOAD;
reg [2:0] INTERNAL_DAC_nLOAD_DONE;
always @ (posedge DAC_REF_CLK) begin
	if(!nRESET) begin
		INTERNAL_DAC_nRESET <= 1'd1;
		INTERNAL_DAC_nRESET_DONE <= 3'b000;
		INTERNAL_DAC_nLOAD <= 1'd1;
		INTERNAL_DAC_nLOAD_DONE <= 3'b000;
	end
	else begin
		if(REG_DAC_CONTROL[1]) begin
			INTERNAL_DAC_nRESET <= 1'd0;
			INTERNAL_DAC_nRESET_DONE <= {INTERNAL_DAC_nRESET_DONE[1:0], 1'd1};
		end
		else begin
			INTERNAL_DAC_nRESET <= 1'd1;
			INTERNAL_DAC_nRESET_DONE <= 3'b000;
		end
		if(REG_DAC_CONTROL[2]) begin
			INTERNAL_DAC_nLOAD <= 1'd0;
			INTERNAL_DAC_nLOAD_DONE <= {INTERNAL_DAC_nLOAD_DONE[1:0] ,1'd1};
		end
		else begin
			INTERNAL_DAC_nLOAD <= 1'd1;
			INTERNAL_DAC_nLOAD_DONE <= 3'b000;
		end
	end
end

assign	DAC_nRST		=	(INTERNAL_DAC_nRESET & nRESET);
assign	DAC_nLOAD	=	(INTERNAL_DAC_nLOAD & EXTERNAL_DAC_nLOAD);

DAC_8734 DAC_8734_inst
(
	.nRESET(nRESET) ,	// input  nRESET_sig
	.DAC_REF_CLK(DAC_REF_CLK) ,	// input  DAC_REF_CLK_sig
	.DAC_SCLK(DAC_SCLK) ,	// output [4:0] DAC_SCLK_sig
	.DAC_nCS(DAC_nCS) ,	// output [4:0] DAC_nCS_sig
	.DAC_SDI(DAC_SDI) ,	// output  DAC_SDI_sig
	.DAC_READY(WIRE_READY) ,	// output  DAC_nREADY_sig
	.DAC_OUTPUT_DONE(WIRE_OUTPUT_DONE) ,	// output  DAC_OUTPUT_DONE_sig
	.DAC_SET_DONE(WIRE_SET_DONE) ,	// output  DAC_SET_DONE_sig
	.REG_DAC_CONTROL(REG_DAC_CONTROL) ,	// input [15:0] REG_DAC_CONTROL_sig
	.REG_DAC0_OUTPUT0(REG_DAC0_OUTPUT0) ,	// input [15:0] REG_DAC0_OUTPUT0_sig
	.REG_DAC0_OUTPUT1(REG_DAC0_OUTPUT1) ,	// input [15:0] REG_DAC0_OUTPUT1_sig
	.REG_DAC0_OUTPUT2(REG_DAC0_OUTPUT2) ,	// input [15:0] REG_DAC0_OUTPUT2_sig
	.REG_DAC0_OUTPUT3(REG_DAC0_OUTPUT3) ,	// input [15:0] REG_DAC0_OUTPUT3_sig
	.REG_DAC1_OUTPUT0(REG_DAC1_OUTPUT0) ,	// input [15:0] REG_DAC1_OUTPUT0_sig
	.REG_DAC1_OUTPUT1(REG_DAC1_OUTPUT1) ,	// input [15:0] REG_DAC1_OUTPUT1_sig
	.REG_DAC1_OUTPUT2(REG_DAC1_OUTPUT2) ,	// input [15:0] REG_DAC1_OUTPUT2_sig
	.REG_DAC1_OUTPUT3(REG_DAC1_OUTPUT3) ,	// input [15:0] REG_DAC1_OUTPUT3_sig
	.REG_DAC2_OUTPUT0(REG_DAC2_OUTPUT0) ,	// input [15:0] REG_DAC2_OUTPUT0_sig
	.REG_DAC2_OUTPUT1(REG_DAC2_OUTPUT1) ,	// input [15:0] REG_DAC2_OUTPUT1_sig
	.REG_DAC2_OUTPUT2(REG_DAC2_OUTPUT2) ,	// input [15:0] REG_DAC2_OUTPUT2_sig
	.REG_DAC2_OUTPUT3(REG_DAC2_OUTPUT3) ,	// input [15:0] REG_DAC2_OUTPUT3_sig
	.REG_DAC3_OUTPUT0(REG_DAC3_OUTPUT0) ,	// input [15:0] REG_DAC3_OUTPUT0_sig
	.REG_DAC3_OUTPUT1(REG_DAC3_OUTPUT1) ,	// input [15:0] REG_DAC3_OUTPUT1_sig
	.REG_DAC3_OUTPUT2(REG_DAC3_OUTPUT2) ,	// input [15:0] REG_DAC3_OUTPUT2_sig
	.REG_DAC3_OUTPUT3(REG_DAC3_OUTPUT3) ,	// input [15:0] REG_DAC3_OUTPUT3_sig
	.REG_DAC4_OUTPUT0(REG_DAC4_OUTPUT0) ,	// input [15:0] REG_DAC4_OUTPUT0_sig
	.REG_DAC4_OUTPUT1(REG_DAC4_OUTPUT1) ,	// input [15:0] REG_DAC4_OUTPUT1_sig
	.REG_DAC4_OUTPUT2(REG_DAC4_OUTPUT2) ,	// input [15:0] REG_DAC4_OUTPUT2_sig
	.REG_DAC4_OUTPUT3(REG_DAC4_OUTPUT3) ,	// input [15:0] REG_DAC4_OUTPUT3_sig
	.REG_DAC_SETCONTROL(REG_DAC_SETCONTROL) ,	// input [15:0] REG_DAC_SETCONTROL_sig
	.REG_DAC_SETBUFFER0(REG_DAC_SETBUFFER0) ,	// input [15:0] REG_DAC_SETBUFFER0_sig
	.REG_DAC_SETBUFFER1(REG_DAC_SETBUFFER1) 	// input [15:0] REG_DAC_SETBUFFER1_sig
);

endmodule
